library verilog;
use verilog.vl_types.all;
entity TB_Clock is
end TB_Clock;
