library verilog;
use verilog.vl_types.all;
entity TB_Parking is
end TB_Parking;
